LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY exception_handler IS PORT(
	input_EXCEPTION_ILLEGAL_INSTRUCTION	: IN STD_LOGIC
); END exception_handler;

ARCHITECTURE gate_level OF exception_handler IS
BEGIN
	-- Deal with exceptions
	
END gate_level;